module hs32_fetch ();
    
endmodule