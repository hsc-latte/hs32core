/**
 * Pipeline Module
 */

module hs32_pipe (
    
);



endmodule