module hs32_reg (

);

endmodule