module top (
    
);
    // Nothing happens here :)
endmodule