module hs32_cpu (
    
);

endmodule
