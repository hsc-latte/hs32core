`include "frontend/sram.v"

module TB_EXT_SRAM();
    
endmodule